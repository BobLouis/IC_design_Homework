library verilog;
use verilog.vl_types.all;
entity testfixture_decoder is
end testfixture_decoder;
