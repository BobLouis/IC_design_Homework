library verilog;
use verilog.vl_types.all;
entity testfixture_encoder is
end testfixture_encoder;
