module LZ77_Encoder(clk,reset,chardata,valid,encode,finish,offset,match_len,char_nxt);

input 				clk;
input 				reset;
input 		[7:0] 	chardata;
output  			valid;
output  			encode;
output  			finish;
output  	[3:0] 	offset;
output  	[2:0] 	match_len;
output  	[7:0] 	char_nxt;

/* write your code here ! */

endmodule
