library verilog;
use verilog.vl_types.all;
entity TB_ELA is
end TB_ELA;
